// sign extend

module sign_extend
(
    input[15:0]     a,
    output[31:0]    out
);
    assign 

endmodule