// i cache
module icache
#(parameter addr_width = 9)
(
	input						nrst,
	input	[addr_width-1:0]	instruction_addr,
	output	[31:0]				instruction_data
);
	reg [31:0] IRAM[2**addr_width-1:0];
	assign instruction_data = IRAM[instruction_addr];
	always @(negedge nrst) begin
		IRAM[0	] = 32'h8c010000;
		IRAM[1	] = 32'h8c020004;
		IRAM[2	] = 32'h8c030008;
		IRAM[3	] = 32'h8c04000c;
		IRAM[4	] = 32'h8c0501f0;
		IRAM[5	] = 32'h8c0601f4;
		IRAM[6	] = 32'h8c0701f8;
		IRAM[7	] = 32'h8c0801fc;
		IRAM[8	] = 32'h00252826;
		IRAM[9	] = 32'h00463026;
		IRAM[10	] = 32'h00673826;
		IRAM[11	] = 32'h00884026;
		IRAM[12	] = 32'h201f0004;
		IRAM[13	] = 32'h20190028;
		IRAM[14	] = 32'h0004dd82;
		IRAM[15	] = 32'h337b03fc;
		IRAM[16	] = 32'h0004e382;
		IRAM[17	] = 32'h339c03fc;
		IRAM[18	] = 32'h0004e982;
		IRAM[19	] = 32'h33bd03fc;
		IRAM[20	] = 32'h8ffa01c4;
		IRAM[21	] = 32'h0004f080;
		IRAM[22	] = 32'h33de03fc;
		IRAM[23	] = 32'h8f9c0200;
		IRAM[24	] = 32'h8fbd0200;
		IRAM[25	] = 32'h8fde0200;
		IRAM[26	] = 32'h8f7b0200;
		IRAM[27	] = 32'h035ce026;
		IRAM[28	] = 32'h001ce600;
		IRAM[29	] = 32'h001dec00;
		IRAM[30	] = 32'h001ef200;
		IRAM[31	] = 32'h039bd820;
		IRAM[32	] = 32'h03bbd820;
		IRAM[33	] = 32'h03dbd820;
		IRAM[34	] = 32'h03610826;
		IRAM[35	] = 32'h00221026;
		IRAM[36	] = 32'h00431826;
		IRAM[37	] = 32'h00642026;
		IRAM[38	] = 32'h00054d82;
		IRAM[39	] = 32'h312903fc;
		IRAM[40	] = 32'h00055382;
		IRAM[41	] = 32'h314a03fc;
		IRAM[42	] = 32'h00055982;
		IRAM[43	] = 32'h316b03fc;
		IRAM[44	] = 32'h00056080;
		IRAM[45	] = 32'h318c03fc;
		IRAM[46	] = 32'h8d290200;
		IRAM[47	] = 32'h8d4a0200;
		IRAM[48	] = 32'h8d6b0200;
		IRAM[49	] = 32'h8d8c0200;
		IRAM[50	] = 32'h00066d82;
		IRAM[51	] = 32'h31ad03fc;
		IRAM[52	] = 32'h00067382;
		IRAM[53	] = 32'h31ce03fc;
		IRAM[54	] = 32'h00067982;
		IRAM[55	] = 32'h31ef03fc;
		IRAM[56	] = 32'h00068080;
		IRAM[57	] = 32'h321003fc;
		IRAM[58	] = 32'h8dad0200;
		IRAM[59	] = 32'h8dce0200;
		IRAM[60	] = 32'h8def0200;
		IRAM[61	] = 32'h8e100200;
		IRAM[62	] = 32'h00078d82;
		IRAM[63	] = 32'h323103fc;
		IRAM[64	] = 32'h00079382;
		IRAM[65	] = 32'h325203fc;
		IRAM[66	] = 32'h00079982;
		IRAM[67	] = 32'h327303fc;
		IRAM[68	] = 32'h0007a080;
		IRAM[69	] = 32'h329403fc;
		IRAM[70	] = 32'h8e310200;
		IRAM[71	] = 32'h8e520200;
		IRAM[72	] = 32'h8e730200;
		IRAM[73	] = 32'h8e940200;
		IRAM[74	] = 32'h0008ad82;
		IRAM[75	] = 32'h32b503fc;
		IRAM[76	] = 32'h0008b382;
		IRAM[77	] = 32'h32d603fc;
		IRAM[78	] = 32'h0008b982;
		IRAM[79	] = 32'h32f703fc;
		IRAM[80	] = 32'h0008c080;
		IRAM[81	] = 32'h331803fc;
		IRAM[82	] = 32'h8eb50200;
		IRAM[83	] = 32'h8ed60200;
		IRAM[84	] = 32'h8ef70200;
		IRAM[85	] = 32'h13f900a0;
		IRAM[86	] = 32'h8f180200;
		IRAM[87	] = 32'h0009d1c2;
		IRAM[88	] = 32'h00092840;
		IRAM[89	] = 32'h101a0002;
		IRAM[90	] = 32'h000ed1c2;
		IRAM[91	] = 32'h38a5011b;
		IRAM[92	] = 32'h000e3040;
		IRAM[93	] = 32'h101a0002;
		IRAM[94	] = 32'h0013d1c2;
		IRAM[95	] = 32'h38c6011b;
		IRAM[96	] = 32'h00133840;
		IRAM[97	] = 32'h101a0002;
		IRAM[98	] = 32'h0018d1c2;
		IRAM[99	] = 32'h38e7011b;
		IRAM[100	] = 32'h00184040;
		IRAM[101	] = 32'h101a0002;
		IRAM[102	] = 32'h00a6d026;
		IRAM[103	] = 32'h3908011b;
		IRAM[104	] = 32'h034ed026;
		IRAM[105	] = 32'h0353d026;
		IRAM[106	] = 32'h0358d026;
		IRAM[107	] = 32'h001ade00;
		IRAM[108	] = 32'h0126d026;
		IRAM[109	] = 32'h0347d026;
		IRAM[110	] = 32'h0353d026;
		IRAM[111	] = 32'h0358d026;
		IRAM[112	] = 32'h001ad400;
		IRAM[113	] = 32'h035bd820;
		IRAM[114	] = 32'h012ed026;
		IRAM[115	] = 32'h0347d026;
		IRAM[116	] = 32'h0348d026;
		IRAM[117	] = 32'h0358d026;
		IRAM[118	] = 32'h001ad200;
		IRAM[119	] = 32'h035bd820;
		IRAM[120	] = 32'h00a9d026;
		IRAM[121	] = 32'h034ed026;
		IRAM[122	] = 32'h0353d026;
		IRAM[123	] = 32'h0348d026;
		IRAM[124	] = 32'h035bd820;
		IRAM[125	] = 32'h000dd1c2;
		IRAM[126	] = 32'h000d2840;
		IRAM[127	] = 32'h101a0002;
		IRAM[128	] = 32'h0012d1c2;
		IRAM[129	] = 32'h38a5011b;
		IRAM[130	] = 32'h00123040;
		IRAM[131	] = 32'h101a0002;
		IRAM[132	] = 32'h0017d1c2;
		IRAM[133	] = 32'h38c6011b;
		IRAM[134	] = 32'h00173840;
		IRAM[135	] = 32'h101a0002;
		IRAM[136	] = 32'h000cd1c2;
		IRAM[137	] = 32'h38e7011b;
		IRAM[138	] = 32'h000c4040;
		IRAM[139	] = 32'h101a0002;
		IRAM[140	] = 32'h00a6d026;
		IRAM[141	] = 32'h3908011b;
		IRAM[142	] = 32'h0352d026;
		IRAM[143	] = 32'h0357d026;
		IRAM[144	] = 32'h034cd026;
		IRAM[145	] = 32'h001ae600;
		IRAM[146	] = 32'h01a6d026;
		IRAM[147	] = 32'h0347d026;
		IRAM[148	] = 32'h0357d026;
		IRAM[149	] = 32'h034cd026;
		IRAM[150	] = 32'h001ad400;
		IRAM[151	] = 32'h035ce020;
		IRAM[152	] = 32'h01b2d026;
		IRAM[153	] = 32'h0347d026;
		IRAM[154	] = 32'h0348d026;
		IRAM[155	] = 32'h034cd026;
		IRAM[156	] = 32'h001ad200;
		IRAM[157	] = 32'h035ce020;
		IRAM[158	] = 32'h00add026;
		IRAM[159	] = 32'h0352d026;
		IRAM[160	] = 32'h0357d026;
		IRAM[161	] = 32'h0348d026;
		IRAM[162	] = 32'h035ce020;
		IRAM[163	] = 32'h0011d1c2;
		IRAM[164	] = 32'h00112840;
		IRAM[165	] = 32'h101a0002;
		IRAM[166	] = 32'h0016d1c2;
		IRAM[167	] = 32'h38a5011b;
		IRAM[168	] = 32'h00163040;
		IRAM[169	] = 32'h101a0002;
		IRAM[170	] = 32'h000bd1c2;
		IRAM[171	] = 32'h38c6011b;
		IRAM[172	] = 32'h000b3840;
		IRAM[173	] = 32'h101a0002;
		IRAM[174	] = 32'h0010d1c2;
		IRAM[175	] = 32'h38e7011b;
		IRAM[176	] = 32'h00104040;
		IRAM[177	] = 32'h101a0002;
		IRAM[178	] = 32'h00a6d026;
		IRAM[179	] = 32'h3908011b;
		IRAM[180	] = 32'h0356d026;
		IRAM[181	] = 32'h034bd026;
		IRAM[182	] = 32'h0350d026;
		IRAM[183	] = 32'h001aee00;
		IRAM[184	] = 32'h0226d026;
		IRAM[185	] = 32'h0347d026;
		IRAM[186	] = 32'h034bd026;
		IRAM[187	] = 32'h0350d026;
		IRAM[188	] = 32'h001ad400;
		IRAM[189	] = 32'h035de820;
		IRAM[190	] = 32'h0236d026;
		IRAM[191	] = 32'h0347d026;
		IRAM[192	] = 32'h0348d026;
		IRAM[193	] = 32'h0350d026;
		IRAM[194	] = 32'h001ad200;
		IRAM[195	] = 32'h035de820;
		IRAM[196	] = 32'h00b1d026;
		IRAM[197	] = 32'h0356d026;
		IRAM[198	] = 32'h034bd026;
		IRAM[199	] = 32'h0348d026;
		IRAM[200	] = 32'h035de820;
		IRAM[201	] = 32'h0015d1c2;
		IRAM[202	] = 32'h00152840;
		IRAM[203	] = 32'h101a0002;
		IRAM[204	] = 32'h000ad1c2;
		IRAM[205	] = 32'h38a5011b;
		IRAM[206	] = 32'h000a3040;
		IRAM[207	] = 32'h101a0002;
		IRAM[208	] = 32'h000fd1c2;
		IRAM[209	] = 32'h38c6011b;
		IRAM[210	] = 32'h000f3840;
		IRAM[211	] = 32'h101a0002;
		IRAM[212	] = 32'h0014d1c2;
		IRAM[213	] = 32'h38e7011b;
		IRAM[214	] = 32'h00144040;
		IRAM[215	] = 32'h101a0002;
		IRAM[216	] = 32'h00a6d026;
		IRAM[217	] = 32'h3908011b;
		IRAM[218	] = 32'h034ad026;
		IRAM[219	] = 32'h034fd026;
		IRAM[220	] = 32'h0354d026;
		IRAM[221	] = 32'h001af600;
		IRAM[222	] = 32'h02a6d026;
		IRAM[223	] = 32'h0347d026;
		IRAM[224	] = 32'h034fd026;
		IRAM[225	] = 32'h0354d026;
		IRAM[226	] = 32'h001ad400;
		IRAM[227	] = 32'h035ef020;
		IRAM[228	] = 32'h02aad026;
		IRAM[229	] = 32'h0347d026;
		IRAM[230	] = 32'h0348d026;
		IRAM[231	] = 32'h0354d026;
		IRAM[232	] = 32'h001ad200;
		IRAM[233	] = 32'h035ef020;
		IRAM[234	] = 32'h00b5d026;
		IRAM[235	] = 32'h034ad026;
		IRAM[236	] = 32'h034fd026;
		IRAM[237	] = 32'h0348d026;
		IRAM[238	] = 32'h035ef020;
		IRAM[239	] = 32'h003b2826;
		IRAM[240	] = 32'h005c3026;
		IRAM[241	] = 32'h007d3826;
		IRAM[242	] = 32'h009e4026;
		IRAM[243	] = 32'h23ff0004;
		IRAM[244	] = 32'h0800000f;
		IRAM[245	] = 32'h0004dd82;
		IRAM[246	] = 32'h00094e00;
		IRAM[247	] = 32'h000e7400;
		IRAM[248	] = 32'h00139a00;
		IRAM[249	] = 32'h012e4820;
		IRAM[250	] = 32'h01334820;
		IRAM[251	] = 32'h01384820;
		IRAM[252	] = 32'h000d6e00;
		IRAM[253	] = 32'h00129400;
		IRAM[254	] = 32'h0017ba00;
		IRAM[255	] = 32'h01b26820;
		IRAM[256	] = 32'h01b76820;
		IRAM[257	] = 32'h01ac6820;
		IRAM[258	] = 32'h00118e00;
		IRAM[259	] = 32'h0016b400;
		IRAM[260	] = 32'h000b5a00;
		IRAM[261	] = 32'h02368820;
		IRAM[262	] = 32'h022b8820;
		IRAM[263	] = 32'h02308820;
		IRAM[264	] = 32'h0015ae00;
		IRAM[265	] = 32'h000a5400;
		IRAM[266	] = 32'h000f7a00;
		IRAM[267	] = 32'h02aaa820;
		IRAM[268	] = 32'h02afa820;
		IRAM[269	] = 32'h02b4a820;
		IRAM[270	] = 32'h00292826;
		IRAM[271	] = 32'h004d3026;
		IRAM[272	] = 32'h00713826;
		IRAM[273	] = 32'h00954026;
		IRAM[274	] = 32'hac050010;
		IRAM[275	] = 32'hac060014;
		IRAM[276	] = 32'hac070018;
		IRAM[277	] = 32'hac08001c;
	end
endmodule
