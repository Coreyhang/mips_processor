module icache(reset,a,rd);
  input reset;
  input[7:0]  a;
  output[31:0]  rd;
  reg[31:0]   RAM[255:0];
  assign rd = RAM[a];
  
  always@(negedge reset)
  begin
    RAM[0  ] = 32'b10001100000001000000000000000000;
	RAM[1  ] = 32'b10001100000001010000000000000001;
	RAM[2  ] = 32'b10001100000001100000000000000010;
	RAM[3  ] = 32'b10001100000001110000000000000011;
	RAM[4  ] = 32'b10001100000100000000000000000100;
	RAM[5  ] = 32'b10001100000100010000000000000101;
	RAM[6  ] = 32'b10001100000100100000000000000110;
	RAM[7  ] = 32'b10001100000100110000000000000111;
	......
	......
	......
  end
  
 
  
endmodule
